package direct_dependency;
endpackage
